class Top#(parameter pckg_sz=32);
mlbx_top_aGENte mlbx_top_aGENte0;


endclass