package Rand_Parameters;
  parameter ROWS = 4;
  parameter COLUMS = 4;
  parameter pckg_sz = 40;
  parameter fifo_depth = 34;
  parameter bdcst = 11111111;
endpackage
