class Top#(parameter pckg_sz=32);

endclass